package shared_pkg;

	logic test_finished;

	// Counters
	integer error_counter=0;
	integer correct_counter=0;

endpackage : shared_pkg